----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    03:11:43 05/22/2022 
-- Design Name: 
-- Module Name:    BRANCH_AND - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity BRANCH_AND is
    Port ( BRANCH_CONTROL : in  STD_LOGIC;
           ZERO : in  STD_LOGIC;
           OUTPUT : out  STD_LOGIC);
end BRANCH_AND;

architecture Behavioral of BRANCH_AND is

begin
OUTPUT <= BRANCH_CONTROL AND ZERO;
end Behavioral;
