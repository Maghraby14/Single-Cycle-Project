----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    03:00:52 05/22/2022 
-- Design Name: 
-- Module Name:    BRANCH_SHIFT_LEFT - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity BRANCH_SHIFT_LEFT is
    Port ( SIGN_EXTEND_OUT : in  STD_LOGIC_VECTOR (31 downto 0);
           OUTPUT : out  STD_LOGIC_VECTOR (31 downto 0));
end BRANCH_SHIFT_LEFT;

architecture Behavioral of BRANCH_SHIFT_LEFT is

begin

OUTPUT <= STD_LOGIC_VECTOR(shift_left(unsigned(SIGN_EXTEND_OUT),2));

end Behavioral;

